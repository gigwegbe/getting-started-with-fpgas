module LED_Toggle_Project
 (input  i_Clk,
  input  i_Switch_1,
  output o_LED_1);
